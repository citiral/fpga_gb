
module system (
	clk_clk,
	reset_reset_n,
	uart_out_rxd,
	uart_out_txd);	

	input		clk_clk;
	input		reset_reset_n;
	input		uart_out_rxd;
	output		uart_out_txd;
endmodule
